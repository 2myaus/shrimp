
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.cpu_types.all;

entity cpu is
end entity;

architecture cpu_a of cpu is
begin

end architecture;

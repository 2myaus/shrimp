library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
package testvec_data is
    constant testvec : std_logic_vector(47 downto 0) := -- 6 bytes
 "100100010001000011111000000000011111111111110000";

end package;
